library ieee;
use ieee.std_logic_1164.all;

package statetype_package is
	type statetype is (s0, s1, s2 ,s3 ,s4 ,s5 ,s6);
end package;

package body statetype_package is
end package body;